magic
tech sky130B
magscale 1 2
timestamp 1662653817
<< obsli1 >>
rect 236104 340159 413848 455521
<< obsm1 >>
rect 1670 3000 582438 703044
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 18 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583432 703610
rect 18 536 583432 703464
rect 18 326 486 536
rect 710 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
rect 165022 326 165994 536
rect 166218 326 167098 536
rect 167322 326 168294 536
rect 168518 326 169490 536
rect 169714 326 170686 536
rect 170910 326 171882 536
rect 172106 326 173078 536
rect 173302 326 174182 536
rect 174406 326 175378 536
rect 175602 326 176574 536
rect 176798 326 177770 536
rect 177994 326 178966 536
rect 179190 326 180162 536
rect 180386 326 181358 536
rect 181582 326 182462 536
rect 182686 326 183658 536
rect 183882 326 184854 536
rect 185078 326 186050 536
rect 186274 326 187246 536
rect 187470 326 188442 536
rect 188666 326 189638 536
rect 189862 326 190742 536
rect 190966 326 191938 536
rect 192162 326 193134 536
rect 193358 326 194330 536
rect 194554 326 195526 536
rect 195750 326 196722 536
rect 196946 326 197826 536
rect 198050 326 199022 536
rect 199246 326 200218 536
rect 200442 326 201414 536
rect 201638 326 202610 536
rect 202834 326 203806 536
rect 204030 326 205002 536
rect 205226 326 206106 536
rect 206330 326 207302 536
rect 207526 326 208498 536
rect 208722 326 209694 536
rect 209918 326 210890 536
rect 211114 326 212086 536
rect 212310 326 213282 536
rect 213506 326 214386 536
rect 214610 326 215582 536
rect 215806 326 216778 536
rect 217002 326 217974 536
rect 218198 326 219170 536
rect 219394 326 220366 536
rect 220590 326 221470 536
rect 221694 326 222666 536
rect 222890 326 223862 536
rect 224086 326 225058 536
rect 225282 326 226254 536
rect 226478 326 227450 536
rect 227674 326 228646 536
rect 228870 326 229750 536
rect 229974 326 230946 536
rect 231170 326 232142 536
rect 232366 326 233338 536
rect 233562 326 234534 536
rect 234758 326 235730 536
rect 235954 326 236926 536
rect 237150 326 238030 536
rect 238254 326 239226 536
rect 239450 326 240422 536
rect 240646 326 241618 536
rect 241842 326 242814 536
rect 243038 326 244010 536
rect 244234 326 245114 536
rect 245338 326 246310 536
rect 246534 326 247506 536
rect 247730 326 248702 536
rect 248926 326 249898 536
rect 250122 326 251094 536
rect 251318 326 252290 536
rect 252514 326 253394 536
rect 253618 326 254590 536
rect 254814 326 255786 536
rect 256010 326 256982 536
rect 257206 326 258178 536
rect 258402 326 259374 536
rect 259598 326 260570 536
rect 260794 326 261674 536
rect 261898 326 262870 536
rect 263094 326 264066 536
rect 264290 326 265262 536
rect 265486 326 266458 536
rect 266682 326 267654 536
rect 267878 326 268758 536
rect 268982 326 269954 536
rect 270178 326 271150 536
rect 271374 326 272346 536
rect 272570 326 273542 536
rect 273766 326 274738 536
rect 274962 326 275934 536
rect 276158 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280626 536
rect 280850 326 281822 536
rect 282046 326 283018 536
rect 283242 326 284214 536
rect 284438 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300682 536
rect 300906 326 301878 536
rect 302102 326 303074 536
rect 303298 326 304270 536
rect 304494 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 308962 536
rect 309186 326 310158 536
rect 310382 326 311354 536
rect 311578 326 312550 536
rect 312774 326 313746 536
rect 313970 326 314942 536
rect 315166 326 316138 536
rect 316362 326 317242 536
rect 317466 326 318438 536
rect 318662 326 319634 536
rect 319858 326 320830 536
rect 321054 326 322026 536
rect 322250 326 323222 536
rect 323446 326 324326 536
rect 324550 326 325522 536
rect 325746 326 326718 536
rect 326942 326 327914 536
rect 328138 326 329110 536
rect 329334 326 330306 536
rect 330530 326 331502 536
rect 331726 326 332606 536
rect 332830 326 333802 536
rect 334026 326 334998 536
rect 335222 326 336194 536
rect 336418 326 337390 536
rect 337614 326 338586 536
rect 338810 326 339782 536
rect 340006 326 340886 536
rect 341110 326 342082 536
rect 342306 326 343278 536
rect 343502 326 344474 536
rect 344698 326 345670 536
rect 345894 326 346866 536
rect 347090 326 347970 536
rect 348194 326 349166 536
rect 349390 326 350362 536
rect 350586 326 351558 536
rect 351782 326 352754 536
rect 352978 326 353950 536
rect 354174 326 355146 536
rect 355370 326 356250 536
rect 356474 326 357446 536
rect 357670 326 358642 536
rect 358866 326 359838 536
rect 360062 326 361034 536
rect 361258 326 362230 536
rect 362454 326 363426 536
rect 363650 326 364530 536
rect 364754 326 365726 536
rect 365950 326 366922 536
rect 367146 326 368118 536
rect 368342 326 369314 536
rect 369538 326 370510 536
rect 370734 326 371614 536
rect 371838 326 372810 536
rect 373034 326 374006 536
rect 374230 326 375202 536
rect 375426 326 376398 536
rect 376622 326 377594 536
rect 377818 326 378790 536
rect 379014 326 379894 536
rect 380118 326 381090 536
rect 381314 326 382286 536
rect 382510 326 383482 536
rect 383706 326 384678 536
rect 384902 326 385874 536
rect 386098 326 387070 536
rect 387294 326 388174 536
rect 388398 326 389370 536
rect 389594 326 390566 536
rect 390790 326 391762 536
rect 391986 326 392958 536
rect 393182 326 394154 536
rect 394378 326 395258 536
rect 395482 326 396454 536
rect 396678 326 397650 536
rect 397874 326 398846 536
rect 399070 326 400042 536
rect 400266 326 401238 536
rect 401462 326 402434 536
rect 402658 326 403538 536
rect 403762 326 404734 536
rect 404958 326 405930 536
rect 406154 326 407126 536
rect 407350 326 408322 536
rect 408546 326 409518 536
rect 409742 326 410714 536
rect 410938 326 411818 536
rect 412042 326 413014 536
rect 413238 326 414210 536
rect 414434 326 415406 536
rect 415630 326 416602 536
rect 416826 326 417798 536
rect 418022 326 418902 536
rect 419126 326 420098 536
rect 420322 326 421294 536
rect 421518 326 422490 536
rect 422714 326 423686 536
rect 423910 326 424882 536
rect 425106 326 426078 536
rect 426302 326 427182 536
rect 427406 326 428378 536
rect 428602 326 429574 536
rect 429798 326 430770 536
rect 430994 326 431966 536
rect 432190 326 433162 536
rect 433386 326 434358 536
rect 434582 326 435462 536
rect 435686 326 436658 536
rect 436882 326 437854 536
rect 438078 326 439050 536
rect 439274 326 440246 536
rect 440470 326 441442 536
rect 441666 326 442546 536
rect 442770 326 443742 536
rect 443966 326 444938 536
rect 445162 326 446134 536
rect 446358 326 447330 536
rect 447554 326 448526 536
rect 448750 326 449722 536
rect 449946 326 450826 536
rect 451050 326 452022 536
rect 452246 326 453218 536
rect 453442 326 454414 536
rect 454638 326 455610 536
rect 455834 326 456806 536
rect 457030 326 458002 536
rect 458226 326 459106 536
rect 459330 326 460302 536
rect 460526 326 461498 536
rect 461722 326 462694 536
rect 462918 326 463890 536
rect 464114 326 465086 536
rect 465310 326 466190 536
rect 466414 326 467386 536
rect 467610 326 468582 536
rect 468806 326 469778 536
rect 470002 326 470974 536
rect 471198 326 472170 536
rect 472394 326 473366 536
rect 473590 326 474470 536
rect 474694 326 475666 536
rect 475890 326 476862 536
rect 477086 326 478058 536
rect 478282 326 479254 536
rect 479478 326 480450 536
rect 480674 326 481646 536
rect 481870 326 482750 536
rect 482974 326 483946 536
rect 484170 326 485142 536
rect 485366 326 486338 536
rect 486562 326 487534 536
rect 487758 326 488730 536
rect 488954 326 489834 536
rect 490058 326 491030 536
rect 491254 326 492226 536
rect 492450 326 493422 536
rect 493646 326 494618 536
rect 494842 326 495814 536
rect 496038 326 497010 536
rect 497234 326 498114 536
rect 498338 326 499310 536
rect 499534 326 500506 536
rect 500730 326 501702 536
rect 501926 326 502898 536
rect 503122 326 504094 536
rect 504318 326 505290 536
rect 505514 326 506394 536
rect 506618 326 507590 536
rect 507814 326 508786 536
rect 509010 326 509982 536
rect 510206 326 511178 536
rect 511402 326 512374 536
rect 512598 326 513478 536
rect 513702 326 514674 536
rect 514898 326 515870 536
rect 516094 326 517066 536
rect 517290 326 518262 536
rect 518486 326 519458 536
rect 519682 326 520654 536
rect 520878 326 521758 536
rect 521982 326 522954 536
rect 523178 326 524150 536
rect 524374 326 525346 536
rect 525570 326 526542 536
rect 526766 326 527738 536
rect 527962 326 528934 536
rect 529158 326 530038 536
rect 530262 326 531234 536
rect 531458 326 532430 536
rect 532654 326 533626 536
rect 533850 326 534822 536
rect 535046 326 536018 536
rect 536242 326 537122 536
rect 537346 326 538318 536
rect 538542 326 539514 536
rect 539738 326 540710 536
rect 540934 326 541906 536
rect 542130 326 543102 536
rect 543326 326 544298 536
rect 544522 326 545402 536
rect 545626 326 546598 536
rect 546822 326 547794 536
rect 548018 326 548990 536
rect 549214 326 550186 536
rect 550410 326 551382 536
rect 551606 326 552578 536
rect 552802 326 553682 536
rect 553906 326 554878 536
rect 555102 326 556074 536
rect 556298 326 557270 536
rect 557494 326 558466 536
rect 558690 326 559662 536
rect 559886 326 560766 536
rect 560990 326 561962 536
rect 562186 326 563158 536
rect 563382 326 564354 536
rect 564578 326 565550 536
rect 565774 326 566746 536
rect 566970 326 567942 536
rect 568166 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572634 536
rect 572858 326 573830 536
rect 574054 326 575026 536
rect 575250 326 576222 536
rect 576446 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580914 536
rect 581138 326 582110 536
rect 582334 326 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 697140 583440 697237
rect 13 697004 583440 697140
rect 13 684484 583586 697004
rect 560 684084 583586 684484
rect 13 684076 583586 684084
rect 13 683676 583440 684076
rect 13 671428 583586 683676
rect 560 671028 583586 671428
rect 13 670884 583586 671028
rect 13 670484 583440 670884
rect 13 658372 583586 670484
rect 560 657972 583586 658372
rect 13 657556 583586 657972
rect 13 657156 583440 657556
rect 13 645316 583586 657156
rect 560 644916 583586 645316
rect 13 644228 583586 644916
rect 13 643828 583440 644228
rect 13 632260 583586 643828
rect 560 631860 583586 632260
rect 13 631036 583586 631860
rect 13 630636 583440 631036
rect 13 619340 583586 630636
rect 560 618940 583586 619340
rect 13 617708 583586 618940
rect 13 617308 583440 617708
rect 13 606284 583586 617308
rect 560 605884 583586 606284
rect 13 604380 583586 605884
rect 13 603980 583440 604380
rect 13 593228 583586 603980
rect 560 592828 583586 593228
rect 13 591188 583586 592828
rect 13 590788 583440 591188
rect 13 580172 583586 590788
rect 560 579772 583586 580172
rect 13 577860 583586 579772
rect 13 577460 583440 577860
rect 13 567116 583586 577460
rect 560 566716 583586 567116
rect 13 564532 583586 566716
rect 13 564132 583440 564532
rect 13 554060 583586 564132
rect 560 553660 583586 554060
rect 13 551340 583586 553660
rect 13 550940 583440 551340
rect 13 541004 583586 550940
rect 560 540604 583586 541004
rect 13 538012 583586 540604
rect 13 537612 583440 538012
rect 13 528084 583586 537612
rect 560 527684 583586 528084
rect 13 524684 583586 527684
rect 13 524284 583440 524684
rect 13 515028 583586 524284
rect 560 514628 583586 515028
rect 13 511492 583586 514628
rect 13 511092 583440 511492
rect 13 501972 583586 511092
rect 560 501572 583586 501972
rect 13 498164 583586 501572
rect 13 497764 583440 498164
rect 13 488916 583586 497764
rect 560 488516 583586 488916
rect 13 484836 583586 488516
rect 13 484436 583440 484836
rect 13 475860 583586 484436
rect 560 475460 583586 475860
rect 13 471644 583586 475460
rect 13 471244 583440 471644
rect 13 462804 583586 471244
rect 560 462404 583586 462804
rect 13 458316 583586 462404
rect 13 457916 583440 458316
rect 13 449748 583586 457916
rect 560 449348 583586 449748
rect 13 444988 583586 449348
rect 13 444588 583440 444988
rect 13 436828 583586 444588
rect 560 436428 583586 436828
rect 13 431796 583586 436428
rect 13 431396 583440 431796
rect 13 423772 583586 431396
rect 560 423372 583586 423772
rect 13 418468 583586 423372
rect 13 418068 583440 418468
rect 13 410716 583586 418068
rect 560 410316 583586 410716
rect 13 405140 583586 410316
rect 13 404740 583440 405140
rect 13 397660 583586 404740
rect 560 397260 583586 397660
rect 13 391948 583586 397260
rect 13 391548 583440 391948
rect 13 384604 583586 391548
rect 560 384204 583586 384604
rect 13 378620 583586 384204
rect 13 378220 583440 378620
rect 13 371548 583586 378220
rect 560 371148 583586 371548
rect 13 365292 583586 371148
rect 13 364892 583440 365292
rect 13 358628 583586 364892
rect 560 358228 583586 358628
rect 13 352100 583586 358228
rect 13 351700 583440 352100
rect 13 345572 583586 351700
rect 560 345172 583586 345572
rect 13 338772 583586 345172
rect 13 338372 583440 338772
rect 13 332516 583586 338372
rect 560 332116 583586 332516
rect 13 325444 583586 332116
rect 13 325044 583440 325444
rect 13 319460 583586 325044
rect 560 319060 583586 319460
rect 13 312252 583586 319060
rect 13 311852 583440 312252
rect 13 306404 583586 311852
rect 560 306004 583586 306404
rect 13 298924 583586 306004
rect 13 298524 583440 298924
rect 13 293348 583586 298524
rect 560 292948 583586 293348
rect 13 285596 583586 292948
rect 13 285196 583440 285596
rect 13 280292 583586 285196
rect 560 279892 583586 280292
rect 13 272404 583586 279892
rect 13 272004 583440 272404
rect 13 267372 583586 272004
rect 560 266972 583586 267372
rect 13 259076 583586 266972
rect 13 258676 583440 259076
rect 13 254316 583586 258676
rect 560 253916 583586 254316
rect 13 245748 583586 253916
rect 13 245348 583440 245748
rect 13 241260 583586 245348
rect 560 240860 583586 241260
rect 13 232556 583586 240860
rect 13 232156 583440 232556
rect 13 228204 583586 232156
rect 560 227804 583586 228204
rect 13 219228 583586 227804
rect 13 218828 583440 219228
rect 13 215148 583586 218828
rect 560 214748 583586 215148
rect 13 205900 583586 214748
rect 13 205500 583440 205900
rect 13 202092 583586 205500
rect 560 201692 583586 202092
rect 13 192708 583586 201692
rect 13 192308 583440 192708
rect 13 189036 583586 192308
rect 560 188636 583586 189036
rect 13 179380 583586 188636
rect 13 178980 583440 179380
rect 13 176116 583586 178980
rect 560 175716 583586 176116
rect 13 166052 583586 175716
rect 13 165652 583440 166052
rect 13 163060 583586 165652
rect 560 162660 583586 163060
rect 13 152860 583586 162660
rect 13 152460 583440 152860
rect 13 150004 583586 152460
rect 560 149604 583586 150004
rect 13 139532 583586 149604
rect 13 139132 583440 139532
rect 13 136948 583586 139132
rect 560 136548 583586 136948
rect 13 126204 583586 136548
rect 13 125804 583440 126204
rect 13 123892 583586 125804
rect 560 123492 583586 123892
rect 13 113012 583586 123492
rect 13 112612 583440 113012
rect 13 110836 583586 112612
rect 560 110436 583586 110836
rect 13 99684 583586 110436
rect 13 99284 583440 99684
rect 13 97780 583586 99284
rect 560 97380 583586 97780
rect 13 86356 583586 97380
rect 13 85956 583440 86356
rect 13 84860 583586 85956
rect 560 84460 583586 84860
rect 13 73164 583586 84460
rect 13 72764 583440 73164
rect 13 71804 583586 72764
rect 560 71404 583586 71804
rect 13 59836 583586 71404
rect 13 59436 583440 59836
rect 13 58748 583586 59436
rect 560 58348 583586 58748
rect 13 46508 583586 58348
rect 13 46108 583440 46508
rect 13 45692 583586 46108
rect 560 45292 583586 45692
rect 13 33316 583586 45292
rect 13 32916 583440 33316
rect 13 32636 583586 32916
rect 560 32236 583586 32636
rect 13 19988 583586 32236
rect 13 19588 583440 19988
rect 13 19580 583586 19588
rect 560 19180 583586 19580
rect 13 6796 583586 19180
rect 13 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583586 6396
rect 13 3299 583586 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 6294 -7654 6914 711590
rect 10794 -7654 11414 711590
rect 15294 -7654 15914 711590
rect 19794 -7654 20414 711590
rect 24294 -7654 24914 711590
rect 28794 -7654 29414 711590
rect 33294 -7654 33914 711590
rect 37794 -7654 38414 711590
rect 42294 -7654 42914 711590
rect 46794 -7654 47414 711590
rect 51294 -7654 51914 711590
rect 55794 -7654 56414 711590
rect 60294 -7654 60914 711590
rect 64794 -7654 65414 711590
rect 69294 -7654 69914 711590
rect 73794 -7654 74414 711590
rect 78294 -7654 78914 711590
rect 82794 -7654 83414 711590
rect 87294 -7654 87914 711590
rect 91794 -7654 92414 711590
rect 96294 -7654 96914 711590
rect 100794 -7654 101414 711590
rect 105294 -7654 105914 711590
rect 109794 -7654 110414 711590
rect 114294 -7654 114914 711590
rect 118794 -7654 119414 711590
rect 123294 -7654 123914 711590
rect 127794 -7654 128414 711590
rect 132294 -7654 132914 711590
rect 136794 -7654 137414 711590
rect 141294 -7654 141914 711590
rect 145794 -7654 146414 711590
rect 150294 -7654 150914 711590
rect 154794 -7654 155414 711590
rect 159294 -7654 159914 711590
rect 163794 -7654 164414 711590
rect 168294 -7654 168914 711590
rect 172794 -7654 173414 711590
rect 177294 -7654 177914 711590
rect 181794 -7654 182414 711590
rect 186294 -7654 186914 711590
rect 190794 -7654 191414 711590
rect 195294 -7654 195914 711590
rect 199794 -7654 200414 711590
rect 204294 -7654 204914 711590
rect 208794 -7654 209414 711590
rect 213294 -7654 213914 711590
rect 217794 -7654 218414 711590
rect 222294 -7654 222914 711590
rect 226794 -7654 227414 711590
rect 231294 -7654 231914 711590
rect 235794 460000 236414 711590
rect 240294 460000 240914 711590
rect 244794 460000 245414 711590
rect 249294 460000 249914 711590
rect 253794 460000 254414 711590
rect 258294 460000 258914 711590
rect 262794 460000 263414 711590
rect 267294 460000 267914 711590
rect 271794 460000 272414 711590
rect 276294 460000 276914 711590
rect 280794 460000 281414 711590
rect 285294 460000 285914 711590
rect 289794 460000 290414 711590
rect 294294 460000 294914 711590
rect 298794 460000 299414 711590
rect 303294 460000 303914 711590
rect 307794 460000 308414 711590
rect 312294 460000 312914 711590
rect 316794 460000 317414 711590
rect 321294 460000 321914 711590
rect 325794 460000 326414 711590
rect 330294 460000 330914 711590
rect 334794 460000 335414 711590
rect 339294 460000 339914 711590
rect 343794 460000 344414 711590
rect 348294 460000 348914 711590
rect 352794 460000 353414 711590
rect 357294 460000 357914 711590
rect 361794 460000 362414 711590
rect 366294 460000 366914 711590
rect 370794 460000 371414 711590
rect 375294 460000 375914 711590
rect 379794 460000 380414 711590
rect 384294 460000 384914 711590
rect 388794 460000 389414 711590
rect 393294 460000 393914 711590
rect 397794 460000 398414 711590
rect 402294 460000 402914 711590
rect 406794 460000 407414 711590
rect 411294 460000 411914 711590
rect 415794 460000 416414 711590
rect 235794 -7654 236414 336000
rect 240294 -7654 240914 336000
rect 244794 -7654 245414 336000
rect 249294 -7654 249914 336000
rect 253794 -7654 254414 336000
rect 258294 -7654 258914 336000
rect 262794 -7654 263414 336000
rect 267294 -7654 267914 336000
rect 271794 -7654 272414 336000
rect 276294 -7654 276914 336000
rect 280794 -7654 281414 336000
rect 285294 -7654 285914 336000
rect 289794 -7654 290414 336000
rect 294294 -7654 294914 336000
rect 298794 -7654 299414 336000
rect 303294 -7654 303914 336000
rect 307794 -7654 308414 336000
rect 312294 -7654 312914 336000
rect 316794 -7654 317414 336000
rect 321294 -7654 321914 336000
rect 325794 -7654 326414 336000
rect 330294 -7654 330914 336000
rect 334794 -7654 335414 336000
rect 339294 -7654 339914 336000
rect 343794 -7654 344414 336000
rect 348294 -7654 348914 336000
rect 352794 -7654 353414 336000
rect 357294 -7654 357914 336000
rect 361794 -7654 362414 336000
rect 366294 -7654 366914 336000
rect 370794 -7654 371414 336000
rect 375294 -7654 375914 336000
rect 379794 -7654 380414 336000
rect 384294 -7654 384914 336000
rect 388794 -7654 389414 336000
rect 393294 -7654 393914 336000
rect 397794 -7654 398414 336000
rect 402294 -7654 402914 336000
rect 406794 -7654 407414 336000
rect 411294 -7654 411914 336000
rect 415794 -7654 416414 336000
rect 420294 -7654 420914 711590
rect 424794 -7654 425414 711590
rect 429294 -7654 429914 711590
rect 433794 -7654 434414 711590
rect 438294 -7654 438914 711590
rect 442794 -7654 443414 711590
rect 447294 -7654 447914 711590
rect 451794 -7654 452414 711590
rect 456294 -7654 456914 711590
rect 460794 -7654 461414 711590
rect 465294 -7654 465914 711590
rect 469794 -7654 470414 711590
rect 474294 -7654 474914 711590
rect 478794 -7654 479414 711590
rect 483294 -7654 483914 711590
rect 487794 -7654 488414 711590
rect 492294 -7654 492914 711590
rect 496794 -7654 497414 711590
rect 501294 -7654 501914 711590
rect 505794 -7654 506414 711590
rect 510294 -7654 510914 711590
rect 514794 -7654 515414 711590
rect 519294 -7654 519914 711590
rect 523794 -7654 524414 711590
rect 528294 -7654 528914 711590
rect 532794 -7654 533414 711590
rect 537294 -7654 537914 711590
rect 541794 -7654 542414 711590
rect 546294 -7654 546914 711590
rect 550794 -7654 551414 711590
rect 555294 -7654 555914 711590
rect 559794 -7654 560414 711590
rect 564294 -7654 564914 711590
rect 568794 -7654 569414 711590
rect 573294 -7654 573914 711590
rect 577794 -7654 578414 711590
rect 582294 -7654 582914 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 228219 3571 231214 461685
rect 231994 459920 235714 461685
rect 236494 459920 240214 461685
rect 240994 459920 244714 461685
rect 245494 459920 249214 461685
rect 249994 459920 253714 461685
rect 254494 459920 258214 461685
rect 258994 459920 262714 461685
rect 263494 459920 267214 461685
rect 267994 459920 271714 461685
rect 272494 459920 276214 461685
rect 276994 459920 280714 461685
rect 281494 459920 285214 461685
rect 285994 459920 289714 461685
rect 290494 459920 294214 461685
rect 294994 459920 298714 461685
rect 299494 459920 303214 461685
rect 303994 459920 307714 461685
rect 308494 459920 312214 461685
rect 312994 459920 316714 461685
rect 317494 459920 321214 461685
rect 321994 459920 325714 461685
rect 326494 459920 330214 461685
rect 330994 459920 334714 461685
rect 335494 459920 339214 461685
rect 339994 459920 343714 461685
rect 344494 459920 348214 461685
rect 348994 459920 352714 461685
rect 353494 459920 357214 461685
rect 357994 459920 361714 461685
rect 362494 459920 366214 461685
rect 366994 459920 370714 461685
rect 371494 459920 375214 461685
rect 375994 459920 379714 461685
rect 380494 459920 384214 461685
rect 384994 459920 388714 461685
rect 389494 459920 393214 461685
rect 393994 459920 397714 461685
rect 398494 459920 402214 461685
rect 402994 459920 406714 461685
rect 407494 459920 411214 461685
rect 411994 459920 415714 461685
rect 416494 459920 420214 461685
rect 231994 336080 420214 459920
rect 231994 3571 235714 336080
rect 236494 3571 240214 336080
rect 240994 3571 244714 336080
rect 245494 3571 249214 336080
rect 249994 3571 253714 336080
rect 254494 3571 258214 336080
rect 258994 3571 262714 336080
rect 263494 3571 267214 336080
rect 267994 3571 271714 336080
rect 272494 3571 276214 336080
rect 276994 3571 280714 336080
rect 281494 3571 285214 336080
rect 285994 3571 289714 336080
rect 290494 3571 294214 336080
rect 294994 3571 298714 336080
rect 299494 3571 303214 336080
rect 303994 3571 307714 336080
rect 308494 3571 312214 336080
rect 312994 3571 316714 336080
rect 317494 3571 321214 336080
rect 321994 3571 325714 336080
rect 326494 3571 330214 336080
rect 330994 3571 334714 336080
rect 335494 3571 339214 336080
rect 339994 3571 343714 336080
rect 344494 3571 348214 336080
rect 348994 3571 352714 336080
rect 353494 3571 357214 336080
rect 357994 3571 361714 336080
rect 362494 3571 366214 336080
rect 366994 3571 370714 336080
rect 371494 3571 375214 336080
rect 375994 3571 379714 336080
rect 380494 3571 384214 336080
rect 384994 3571 388714 336080
rect 389494 3571 393214 336080
rect 393994 3571 397714 336080
rect 398494 3571 402214 336080
rect 402994 3571 406714 336080
rect 407494 3571 411214 336080
rect 411994 3571 415714 336080
rect 416494 3571 420214 336080
rect 420994 3571 423693 461685
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 700366 592650 700986
rect -8726 695866 592650 696486
rect -8726 691366 592650 691986
rect -8726 686866 592650 687486
rect -8726 682366 592650 682986
rect -8726 677866 592650 678486
rect -8726 673366 592650 673986
rect -8726 668866 592650 669486
rect -8726 664366 592650 664986
rect -8726 659866 592650 660486
rect -8726 655366 592650 655986
rect -8726 650866 592650 651486
rect -8726 646366 592650 646986
rect -8726 641866 592650 642486
rect -8726 637366 592650 637986
rect -8726 632866 592650 633486
rect -8726 628366 592650 628986
rect -8726 623866 592650 624486
rect -8726 619366 592650 619986
rect -8726 614866 592650 615486
rect -8726 610366 592650 610986
rect -8726 605866 592650 606486
rect -8726 601366 592650 601986
rect -8726 596866 592650 597486
rect -8726 592366 592650 592986
rect -8726 587866 592650 588486
rect -8726 583366 592650 583986
rect -8726 578866 592650 579486
rect -8726 574366 592650 574986
rect -8726 569866 592650 570486
rect -8726 565366 592650 565986
rect -8726 560866 592650 561486
rect -8726 556366 592650 556986
rect -8726 551866 592650 552486
rect -8726 547366 592650 547986
rect -8726 542866 592650 543486
rect -8726 538366 592650 538986
rect -8726 533866 592650 534486
rect -8726 529366 592650 529986
rect -8726 524866 592650 525486
rect -8726 520366 592650 520986
rect -8726 515866 592650 516486
rect -8726 511366 592650 511986
rect -8726 506866 592650 507486
rect -8726 502366 592650 502986
rect -8726 497866 592650 498486
rect -8726 493366 592650 493986
rect -8726 488866 592650 489486
rect -8726 484366 592650 484986
rect -8726 479866 592650 480486
rect -8726 475366 592650 475986
rect -8726 470866 592650 471486
rect -8726 466366 592650 466986
rect -8726 461866 592650 462486
rect -8726 457366 592650 457986
rect -8726 452866 592650 453486
rect -8726 448366 592650 448986
rect -8726 443866 592650 444486
rect -8726 439366 592650 439986
rect -8726 434866 592650 435486
rect -8726 430366 592650 430986
rect -8726 425866 592650 426486
rect -8726 421366 592650 421986
rect -8726 416866 592650 417486
rect -8726 412366 592650 412986
rect -8726 407866 592650 408486
rect -8726 403366 592650 403986
rect -8726 398866 592650 399486
rect -8726 394366 592650 394986
rect -8726 389866 592650 390486
rect -8726 385366 592650 385986
rect -8726 380866 592650 381486
rect -8726 376366 592650 376986
rect -8726 371866 592650 372486
rect -8726 367366 592650 367986
rect -8726 362866 592650 363486
rect -8726 358366 592650 358986
rect -8726 353866 592650 354486
rect -8726 349366 592650 349986
rect -8726 344866 592650 345486
rect -8726 340366 592650 340986
rect -8726 335866 592650 336486
rect -8726 331366 592650 331986
rect -8726 326866 592650 327486
rect -8726 322366 592650 322986
rect -8726 317866 592650 318486
rect -8726 313366 592650 313986
rect -8726 308866 592650 309486
rect -8726 304366 592650 304986
rect -8726 299866 592650 300486
rect -8726 295366 592650 295986
rect -8726 290866 592650 291486
rect -8726 286366 592650 286986
rect -8726 281866 592650 282486
rect -8726 277366 592650 277986
rect -8726 272866 592650 273486
rect -8726 268366 592650 268986
rect -8726 263866 592650 264486
rect -8726 259366 592650 259986
rect -8726 254866 592650 255486
rect -8726 250366 592650 250986
rect -8726 245866 592650 246486
rect -8726 241366 592650 241986
rect -8726 236866 592650 237486
rect -8726 232366 592650 232986
rect -8726 227866 592650 228486
rect -8726 223366 592650 223986
rect -8726 218866 592650 219486
rect -8726 214366 592650 214986
rect -8726 209866 592650 210486
rect -8726 205366 592650 205986
rect -8726 200866 592650 201486
rect -8726 196366 592650 196986
rect -8726 191866 592650 192486
rect -8726 187366 592650 187986
rect -8726 182866 592650 183486
rect -8726 178366 592650 178986
rect -8726 173866 592650 174486
rect -8726 169366 592650 169986
rect -8726 164866 592650 165486
rect -8726 160366 592650 160986
rect -8726 155866 592650 156486
rect -8726 151366 592650 151986
rect -8726 146866 592650 147486
rect -8726 142366 592650 142986
rect -8726 137866 592650 138486
rect -8726 133366 592650 133986
rect -8726 128866 592650 129486
rect -8726 124366 592650 124986
rect -8726 119866 592650 120486
rect -8726 115366 592650 115986
rect -8726 110866 592650 111486
rect -8726 106366 592650 106986
rect -8726 101866 592650 102486
rect -8726 97366 592650 97986
rect -8726 92866 592650 93486
rect -8726 88366 592650 88986
rect -8726 83866 592650 84486
rect -8726 79366 592650 79986
rect -8726 74866 592650 75486
rect -8726 70366 592650 70986
rect -8726 65866 592650 66486
rect -8726 61366 592650 61986
rect -8726 56866 592650 57486
rect -8726 52366 592650 52986
rect -8726 47866 592650 48486
rect -8726 43366 592650 43986
rect -8726 38866 592650 39486
rect -8726 34366 592650 34986
rect -8726 29866 592650 30486
rect -8726 25366 592650 25986
rect -8726 20866 592650 21486
rect -8726 16366 592650 16986
rect -8726 11866 592650 12486
rect -8726 7366 592650 7986
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 336000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 460000 254414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 336000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 460000 290414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 336000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 460000 326414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 336000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 460000 362414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 336000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 460000 398414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 336000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 262794 460000 263414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 336000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 298794 460000 299414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 336000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 334794 460000 335414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 336000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 370794 460000 371414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 336000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 406794 460000 407414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 235794 460000 236414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 271794 460000 272414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 307794 460000 308414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 343794 460000 344414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 379794 460000 380414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 336000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 415794 460000 416414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 336000 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 244794 460000 245414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 336000 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 280794 460000 281414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 336000 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 316794 460000 317414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 336000 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 352794 460000 353414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 336000 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 388794 460000 389414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 336000 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 240294 460000 240914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 336000 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 276294 460000 276914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 336000 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 312294 460000 312914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 336000 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 348294 460000 348914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 336000 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 384294 460000 384914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 336000 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 249294 460000 249914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 336000 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 285294 460000 285914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 336000 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 321294 460000 321914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 336000 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 357294 460000 357914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 336000 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 393294 460000 393914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 336000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 258294 460000 258914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 336000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 294294 460000 294914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 336000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 330294 460000 330914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 336000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 366294 460000 366914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 336000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 402294 460000 402914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 336000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 267294 460000 267914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 336000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 303294 460000 303914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 336000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 339294 460000 339914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 336000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 375294 460000 375914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 336000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 411294 460000 411914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9683374
string GDS_FILE /home/nvm_user4/usr/mpw_7_files/caravel_user_project_analog/openlane/user_analog_project_wrapper/runs/22_09_08_21_44/results/signoff/user_analog_project_wrapper.magic.gds
string GDS_START 7854180
<< end >>

